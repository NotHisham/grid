// =================================================================================
// Verilog Code for an Electric Vehicle (EV) Charging System
//
// ADVANCED VERSION: This code uses more complex cryptographic functions.
// INCLUDES TIMESTAMPS: Incorporates timestamps and time-lag checks to prevent replay attacks.
// FLOWCHART ALIGNED: Logic and variable names updated to match the provided flowcharts.
//
// The code is split into three modules:
// 1. EV Registration
// 2. CS Registration
// 3. EV-CS Authentication
// =================================================================================


// =================================================================================
// MODULE 1: EV Registration with the Utility Service Provider (USP)
// This module follows "Table 1: Registration of EV with USP" from the flowchart.
// =================================================================================
module EV_USP_Registration (
    input clk,                  /* Clock signal to synchronize operations */
    input rst,                  /* Reset signal to clear all values */
    input [63:0] ev_id_i,       /* Input: The EV's unique, real Identity (IDi) */
    input [63:0] ev_ch_i,       /* Input: The EV's secret Challenge value (CHi), which acts as a nonce. */
    input [63:0] usp_pub_key_j, /* Input: The USP's Public Key, used for encryption */
    input [63:0] T1,            /* Input: The EV's timestamp (T1) for the initial message */
    output reg [255:0] M1,      /* Output: The first message (PSIDEVi, CHi, RSi, T1) sent from the EV to the USP */
    output reg [255:0] M2,      /* Output: The second message (Aj, IDj, Pubj, T2) sent back from the USP to the EV */
    output reg registration_complete, /* A flag that goes high when done */
    output reg registration_failed    /* A flag that goes high if the timestamp check fails */
);

    /* --- Parameters --- */
    parameter ACCEPTABLE_DELAY = 10; /* Max allowed time units (delta t) between message send and receive */

    /* Internal wires and registers to hold intermediate values during the process. */
    reg [63:0] rs_i;
    reg [63:0] psidev_i;
    reg [63:0] a_j;
    reg [63:0] usp_id_j;
    reg [63:0] decrypted_aj;
    reg [63:0] decrypted_idj;
    reg [63:0] decrypted_pubj;
    reg [63:0] received_t1;
    reg [63:0] received_t2;
    reg [63:0] T2; // Timestamp generated by USP
    reg [63:0] TS2; // Timestamp at USP when M1 is received
    reg [63:0] TS3; // Timestamp at EV when M2 is received
    
    // Temporary registers to hold full decrypted message before unpacking
    reg [255:0] temp_m1_decrypted;
    reg [255:0] temp_m2_decrypted;


    /* An advanced model of a Physically Unclonable Function (PUF) */
    function [63:0] puf (input [63:0] challenge);
        reg [63:0] lfsr_reg; integer i;
        begin
            lfsr_reg = challenge;
            for (i = 0; i < 64; i = i + 1) begin
                lfsr_reg = {lfsr_reg[62:0], lfsr_reg[63] ^ lfsr_reg[62] ^ lfsr_reg[60] ^ lfsr_reg[59]};
            end
            puf = lfsr_reg;
        end
    endfunction

    /* An advanced model of a Hash function. Now takes 320 bits to include Pubj */
    function [63:0] hash (input [319:0] data);
        reg [63:0] state; reg [63:0] round_key; integer i; reg [63:0] data_chunk;
        begin
            state = 64'hA5A5A5A5A5A5A5A5;
            for (i = 0; i < 5; i = i + 1) begin
                case(i)
                    0: data_chunk = data[63:0]; 1: data_chunk = data[127:64]; 2: data_chunk = data[191:128];
                    3: data_chunk = data[255:192]; 4: data_chunk = data[319:256];
                    default: data_chunk = 64'h0;
                endcase
                state = state ^ data_chunk;
                round_key = 64'hC3C3C3C3C3C3C3C3 >> (i * 7);
                state = (state <<< 3) ^ (state >> 5) ^ round_key;
            end
            hash = state;
        end
    endfunction
    
    /* Encryption/Decryption model using XOR, size updated to 256 bits for M1 and M2. */
    function [255:0] encrypt (input [255:0] plaintext, input [63:0] key);
        encrypt = plaintext ^ {4{key}};
    endfunction

    always @(posedge clk or posedge rst) begin
        if (rst) begin
            M1 <= 0; M2 <= 0; registration_complete <= 0; registration_failed <= 0;
            rs_i <= 0; psidev_i <= 0; a_j <= 0;
        end else begin
            /* === EV SIDE: Step 1 - Preparation === */
            rs_i <= puf(ev_ch_i);
            psidev_i <= hash({ev_id_i, rs_i, 192'd0}); // Pad to 320 bits for hash function
            M1 <= encrypt({psidev_i, ev_ch_i, rs_i, T1}, usp_pub_key_j);

            /* === USP SIDE: Step 2 - Verification and Response === */
            /* USP decrypts M1 to get the contents and the timestamp T1 */
            temp_m1_decrypted = encrypt(M1, usp_pub_key_j);
            received_t1 = temp_m1_decrypted[63:0];
            
            /* USP checks if the message is recent. TS2 is the USP's current time. */
            TS2 <= T1 + 5; // Simulating network delay
            
            if ((TS2 - received_t1) > ACCEPTABLE_DELAY) begin
                registration_failed <= 1;
                registration_complete <= 0;
            end else begin
                registration_failed <= 0;
                
                /* Timestamp is valid, so USP proceeds. */
                usp_id_j <= 64'hABCDEF9876543210;
                /* Aj = H(IDi || CHi || RSi || IDj || Pubj) as per flowchart */
                a_j <= hash({ev_id_i, ev_ch_i, rs_i, usp_id_j, usp_pub_key_j});

                /* USP generates its own timestamp, T2, for the response message. */
                T2 <= TS2 + 1;

                /* USP sends M2 = E(Aj, IDj, Pubj, T2) using EV's public key (IDi for this simple model) */
                M2 <= encrypt({a_j, usp_id_j, usp_pub_key_j, T2}, ev_id_i);

                /* === EV SIDE: Step 3 - Finalization === */
                /* EV decrypts M2 to get the contents and the timestamp T2 */
                temp_m2_decrypted = encrypt(M2, ev_id_i);
                {decrypted_aj, decrypted_idj, decrypted_pubj, received_t2} = temp_m2_decrypted;

                /* EV checks if the USP's response is recent. TS3 is the EV's current time. */
                TS3 <= T2 + 6; // Simulating another small network delay

                if ((TS3 - received_t2) > ACCEPTABLE_DELAY) begin
                    registration_failed <= 1;
                    registration_complete <= 0;
                end else begin
                    /* Timestamp is valid, registration is successful. */
                    registration_failed <= 0;
                    registration_complete <= 1;
                end
            end
        end
    end
endmodule


// =================================================================================
// MODULE 2: CS Registration with the Utility Service Provider (USP)
// This module follows "Table 2: Registration of CS with USP" from the flowchart.
// =================================================================================
module CS_USP_Registration (
    input clk,
    input rst,
    input [63:0] cs_id_k,
    input [63:0] cs_ch_k,       /* Input: The CS's secret Challenge value (CHk), which acts as a nonce. */
    input [63:0] cs_rs_k,
    input [63:0] cs_pub_key_k,
    input [63:0] usp_pub_key_j,
    input [63:0] T1,         /* Input: The CS's timestamp (T1) for the initial message */
    output reg [319:0] M1,   /* Output: Message 1 (IDk, CHk, RSk, Pubk, T1) */
    output reg [191:0] M2,   /* Output: Message 2 (IDj, Aj, T2) */
    output reg registration_complete,
    output reg registration_failed
);
    
    parameter ACCEPTABLE_DELAY = 10;
    reg [63:0] a_j;
    reg [63:0] usp_id_j;
    reg [63:0] decrypted_aj;
    reg [63:0] decrypted_idj;
    reg [63:0] received_t1;
    reg [63:0] received_t2;
    reg [63:0] T2;
    reg [63:0] TS2; // Timestamp at USP
    reg [63:0] TS3; // Timestamp at CS
    
    // Temporary registers to hold full decrypted message before unpacking
    reg [319:0] temp_m1_decrypted;
    reg [191:0] temp_m2_decrypted;

    /* Hash function for 384-bit input to include all terms for Aj */
    function [63:0] hash (input [383:0] data);
        reg [63:0] state; reg [63:0] round_key; integer i; reg [63:0] data_chunk;
        begin
            state = 64'hA5A5A5A5A5A5A5A5;
            for (i = 0; i < 6; i = i + 1) begin
                case(i)
                    0: data_chunk = data[63:0]; 1: data_chunk = data[127:64]; 2: data_chunk = data[191:128];
                    3: data_chunk = data[255:192]; 4: data_chunk = data[319:256]; 5: data_chunk = data[383:320];
                    default: data_chunk = 64'h0;
                endcase
                state = state ^ data_chunk;
                round_key = 64'hC3C3C3C3C3C3C3C3 >> (i * 6);
                state = (state <<< 3) ^ (state >> 5) ^ round_key;
            end
            hash = state;
        end
    endfunction

    function [319:0] encrypt_m1 (input [319:0] plaintext, input [63:0] key);
        encrypt_m1 = plaintext ^ {5{key}};
    endfunction
    function [191:0] encrypt_m2 (input [191:0] plaintext, input [63:0] key);
        encrypt_m2 = plaintext ^ {3{key}};
    endfunction

    always @(posedge clk or posedge rst) begin
        if (rst) begin
            M1 <= 0; M2 <= 0; registration_complete <= 0; registration_failed <= 0; a_j <= 0; usp_id_j <= 0;
        end else begin
            /* === CS SIDE: Step 1 - Preparation === */
            M1 <= encrypt_m1({cs_id_k, cs_ch_k, cs_rs_k, cs_pub_key_k, T1}, usp_pub_key_j);

            /* === USP SIDE: Step 2 - Verification and Response === */
            temp_m1_decrypted = encrypt_m1(M1, usp_pub_key_j);
            received_t1 = temp_m1_decrypted[63:0];
            TS2 <= T1 + 4; // Simulating network delay

            if ((TS2 - received_t1) > ACCEPTABLE_DELAY) begin
                registration_failed <= 1;
                registration_complete <= 0;
            end else begin
                registration_failed <= 0;
                usp_id_j <= 64'hFEDCBA0987654321;
                /* Aj = H(IDk || CHk || RSk || IDj || Pubj || Pubk) as per flowchart */
                a_j <= hash({cs_id_k, cs_ch_k, cs_rs_k, usp_id_j, usp_pub_key_j, cs_pub_key_k});
                T2 <= TS2 + 1;
                M2 <= encrypt_m2({usp_id_j, a_j, T2}, cs_pub_key_k);

                /* === CS SIDE: Step 3 - Finalization === */
                temp_m2_decrypted = encrypt_m2(M2, cs_pub_key_k);
                {decrypted_idj, decrypted_aj, received_t2} = temp_m2_decrypted;
                TS3 <= T2 + 5; // Simulating return network delay
                
                if ((TS3 - received_t2) > ACCEPTABLE_DELAY) begin
                    registration_failed <= 1;
                    registration_complete <= 0;
                end else begin
                    registration_failed <= 0;
                    registration_complete <= 1;
                end
            end
        end
    end
endmodule

// =================================================================================
// MODULE 3: EV-CS Authentication
// This module follows "Table 2: Authentication between EV and CS" from the flowchart.
// =================================================================================
module EV_CS_Authentication (
    input clk,
    input rst,
    input [63:0] ev_psidev_i,
    input [63:0] ev_pub_key,
    input [63:0] cs_pub_key,
    input [63:0] ev_retrieved_rs_i,
    output reg mutual_authentication_established,
    output reg authentication_failed
);
    
    parameter ACCEPTABLE_DELAY = 10;

    reg [63:0] ev_n1, cs_n2, cs_n4;
    reg [63:0] T1, T2, T3, T4;
    reg [63:0] TS2, TS3, TS4, TS5; // Timestamps at point of reception
    
    /* Messages exchanged between EV and CS, sizes updated to match flowchart */
    reg [255:0] m1; reg [319:0] m2; reg [383:0] m3; reg [447:0] m4;
    
    reg [63:0] cs_ch_k, cs_seed, cs_k_k, cs_id_k, token_tk_k, rs_k_prime, k_sk;
    wire [63:0] ev_ch_k; // This is the challenge (nonce) from the CS
    reg [63:0] ev_ka; // Renamed from ev_k_i to match flowchart
    reg [63:0] received_rsk;
    reg ev_cs_verified;
    
    reg t1_valid, t2_valid, t3_valid, t4_valid;
    
    // Temporary registers to hold full decrypted messages before unpacking
    reg [255:0] temp_m1_decrypted_auth;
    reg [319:0] temp_m2_decrypted_auth;
    reg [383:0] temp_m3_decrypted_auth;
    reg [447:0] temp_m4_decrypted_auth;

    function [63:0] puf (input [63:0] challenge);
        reg [63:0] lfsr_reg; integer i;
        begin lfsr_reg = challenge; for (i = 0; i < 64; i = i + 1) lfsr_reg = {lfsr_reg[62:0], lfsr_reg[63] ^ lfsr_reg[62] ^ lfsr_reg[60] ^ lfsr_reg[59]}; puf = lfsr_reg; end
    endfunction

    function [63:0] hash (input [191:0] data);
        reg [63:0] state; reg [63:0] round_key; integer i; reg [63:0] data_chunk;
        begin state = 64'hA5A5A5A5A5A5A5A5; for (i = 0; i < 3; i = i + 1) begin case(i) 0: data_chunk = data[63:0]; 1: data_chunk = data[127:64]; 2: data_chunk = data[191:128]; default: data_chunk = 64'h0; endcase state = state ^ data_chunk; round_key = 64'hC3C3C3C3C3C3C3C3 >> (i * 9); state = (state <<< 3) ^ (state >> 5) ^ round_key; end hash = state; end
    endfunction

    /* Encryption functions with updated sizes */
    function [255:0] encrypt_m1 (input [255:0] plaintext, input [63:0] key); encrypt_m1 = plaintext ^ {4{key}}; endfunction
    function [319:0] encrypt_m2 (input [319:0] plaintext, input [63:0] key); encrypt_m2 = plaintext ^ {5{key}}; endfunction
    function [383:0] encrypt_m3 (input [383:0] plaintext, input [63:0] key); encrypt_m3 = plaintext ^ {6{key}}; endfunction
    function [447:0] encrypt_m4 (input [447:0] plaintext, input [63:0] key); encrypt_m4 = plaintext ^ {7{key}}; endfunction

    /* Continuous assignments for extracting values from decrypted messages */
    wire [319:0] temp_m2_decrypted_wire;
    assign temp_m2_decrypted_wire = encrypt_m2(m2, ev_pub_key);
    assign ev_ch_k = temp_m2_decrypted_wire[255:192]; // Position of CHk in M2

    always @(posedge clk or posedge rst) begin
        if (rst) begin
            mutual_authentication_established <= 0; authentication_failed <= 0; ev_ka <= 0; ev_cs_verified <= 0;
            t1_valid <= 0; t2_valid <= 0; t3_valid <= 0; t4_valid <= 0;
        end else begin
            /* === STEP 1: EV sends M1 to CS === */
            ev_n1 <= 64'h1111_1111_1111_1111;
            T1 <= 100; // EV sends message at time 100
            m1 <= encrypt_m1({ev_psidev_i, ev_n1, ev_pub_key, T1}, cs_pub_key);

            /* --- CS receives M1 and checks timestamp T1 --- */
            reg [63:0] received_t1;
            TS2 = T1 + 5; // Simulate current time at CS
            temp_m1_decrypted_auth = encrypt_m1(m1, cs_pub_key);
            received_t1 = temp_m1_decrypted_auth[63:0];
            t1_valid <= ((TS2 - received_t1) <= ACCEPTABLE_DELAY);
            
            if (!t1_valid) begin authentication_failed <= 1;
            end else begin
                /* === STEP 2: CS sends back M2 === */
                cs_ch_k <= 64'hAAAAAAAAAAAAAAAA; // This challenge (nonce) should be random in a real implementation.
                cs_seed <= 64'hBBBBBBBBBBBBBBBB;
                cs_n2   <= 64'h2222_2222_2222_2222;
                cs_id_k <= 64'hDDDDDDDDDDDDDDDD;
                T2 <= TS2 + 1;
                m2 <= encrypt_m2({cs_id_k, cs_ch_k, cs_n2, cs_seed, T2}, ev_pub_key);

                /* --- EV receives M2 and checks timestamp T2 --- */
                reg [63:0] received_t2;
                TS3 = T2 + 4; // Simulate current time at EV
                temp_m2_decrypted_auth = encrypt_m2(m2, ev_pub_key);
                received_t2 = temp_m2_decrypted_auth[63:0];
                t2_valid <= ((TS3 - received_t2) <= ACCEPTABLE_DELAY);

                if (!t2_valid) begin authentication_failed <= 1;
                end else begin
                    /* === STEP 3: EV sends M3 === */
                    reg [63:0] seed_from_m2;
                    seed_from_m2 = temp_m2_decrypted_auth[127:64];
                    ev_ka <= puf(seed_from_m2); // Ka = PUF(seed) as per flowchart
                    T3 <= TS3 + 1;
                    /* M3 = E(PSIDEVi, N1, RSi, CHk, Ka, T3)Pubk */
                    m3 <= encrypt_m3({ev_psidev_i, ev_n1, ev_retrieved_rs_i, ev_ch_k, ev_ka, T3}, cs_pub_key);

                    /* --- CS receives M3 and checks timestamp T3 --- */
                    reg [63:0] received_t3;
                    TS4 = T3 + 6; // Simulate current time at CS
                    temp_m3_decrypted_auth = encrypt_m3(m3, cs_pub_key);
                    received_t3 = temp_m3_decrypted_auth[63:0];
                    t3_valid <= ((TS4 - received_t3) <= ACCEPTABLE_DELAY);

                    if (!t3_valid) begin authentication_failed <= 1;
                    end else begin
                        /* === STEP 4: CS authenticates EV and sends final message M4 === */
                        token_tk_k <= hash({ev_psidev_i, ev_retrieved_rs_i, cs_id_k});
                        rs_k_prime <= puf(cs_ch_k); // This is RSk
                        cs_k_k <= puf(cs_seed);
                        k_sk <= hash({cs_k_k, 128'd0}); // This is Ksk
                        cs_n4 <= 64'h4444_4444_4444_4444;
                        T4 <= TS4 + 1;
                        /* M4 = E(IDk, CHk, N4, RSk, TKk, Ksk, T4)Ka */
                        m4 <= encrypt_m4({cs_id_k, cs_ch_k, cs_n4, rs_k_prime, token_tk_k, k_sk, T4}, ev_ka);
                        
                        /* --- EV receives M4 and checks timestamp T4 --- */
                        reg [63:0] received_t4;
                        TS5 = T4 + 5;
                        temp_m4_decrypted_auth = encrypt_m4(m4, ev_ka);
                        received_t4 = temp_m4_decrypted_auth[63:0];
                        t4_valid <= ((TS5 - received_t4) <= ACCEPTABLE_DELAY);
                        
                        if (!t4_valid) begin authentication_failed <= 1;
                        end else begin
                           /* === FINAL STEP: EV verifies CS's final response by checking RSk === */
                           received_rsk = temp_m4_decrypted_auth[255:192];
                           
                           if (received_rsk == puf(ev_ch_k)) begin
                               ev_cs_verified <= 1;
                               mutual_authentication_established <= 1;
                               authentication_failed <= 0;
                           end else begin
                               ev_cs_verified <= 0;
                               mutual_authentication_established <= 0;
                               authentication_failed <= 1;
                           end
                        end
                    end
                end
            end
        end
    end
endmodule
